hihi

im testing something not important
