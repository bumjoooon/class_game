hihi

iam testing something not important




what am i doing now?

this work done in untracked file
this work done in tracked file

add this line after reset hard
