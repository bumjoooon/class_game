hihi

iam testing something not important


what am i doing now?


add this line after reset hard
