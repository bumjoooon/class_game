hihi

iam testing something not important


what am i doing now?
